// This is the unpowered netlist.
module top (clk,
    convst_bar,
    duty_high,
    duty_low,
    rst,
    data_in);
 input clk;
 output convst_bar;
 output duty_high;
 output duty_low;
 input rst;
 input [7:0] data_in;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire \clkdivider.clk2[0] ;
 wire \clkdivider.clk2[1] ;
 wire \clkdivider.clk2[2] ;
 wire \clkdivider.clk2[3] ;
 wire \clkdivider.clk2[4] ;
 wire \clkdivider.clk2[5] ;
 wire \clkdivider.clk_comp ;
 wire \clkdivider.clk_dpwm ;
 wire \clkdivider.count[0] ;
 wire \clkdivider.count[1] ;
 wire \clkdivider.count[2] ;
 wire \clkdivider.count[3] ;
 wire \clkdivider.count[4] ;
 wire \clkdivider.count[5] ;
 wire \clkdivider.count[6] ;
 wire clknet_0_clk;
 wire clknet_1_0__leaf_clk;
 wire clknet_1_1__leaf_clk;
 wire \dither.count[0] ;
 wire \dither.count[1] ;
 wire \dither.count[2] ;
 wire \dither.d_n_input[0] ;
 wire \dither.d_n_input[1] ;
 wire \dither.d_n_input[2] ;
 wire \dither.d_n_input[3] ;
 wire \dither.d_n_input[4] ;
 wire \dither.d_n_input[5] ;
 wire \dither.d_n_input[6] ;
 wire \dither.d_n_input[7] ;
 wire \dither.d_n_input[8] ;
 wire \encoder.en[0] ;
 wire \encoder.en[1] ;
 wire \encoder.en[2] ;
 wire \encoder.en[3] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \stanley.d_n_1[0] ;
 wire \stanley.d_n_1[10] ;
 wire \stanley.d_n_1[11] ;
 wire \stanley.d_n_1[12] ;
 wire \stanley.d_n_1[13] ;
 wire \stanley.d_n_1[14] ;
 wire \stanley.d_n_1[15] ;
 wire \stanley.d_n_1[1] ;
 wire \stanley.d_n_1[2] ;
 wire \stanley.d_n_1[3] ;
 wire \stanley.d_n_1[4] ;
 wire \stanley.d_n_1[5] ;
 wire \stanley.d_n_1[6] ;
 wire \stanley.d_n_1[7] ;
 wire \stanley.d_n_1[8] ;
 wire \stanley.d_n_1[9] ;
 wire \stanley.d_n_reg[0] ;
 wire \stanley.d_n_reg[1] ;
 wire \stanley.d_n_reg[2] ;
 wire \stanley.d_n_reg[3] ;
 wire \stanley.d_n_reg[4] ;
 wire \stanley.d_n_reg[5] ;
 wire \stanley.en1[0] ;
 wire \stanley.en1[1] ;
 wire \stanley.en1[2] ;
 wire \stanley.en1[3] ;
 wire \stanley.en2[0] ;
 wire \stanley.en2[1] ;
 wire \stanley.en2[2] ;
 wire \stanley.en2[3] ;
 wire \stanley.en3[0] ;
 wire \stanley.en3[1] ;
 wire \stanley.en3[2] ;
 wire \stanley.en3[3] ;
 wire \stanley.en[0] ;
 wire \stanley.en[1] ;
 wire \stanley.en[2] ;
 wire \stanley.en[3] ;

 sky130_fd_sc_hd__decap_8 FILLER_0_0_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_90 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__and3_1 _0550_ (.A(\clkdivider.clk2[1] ),
    .B(\clkdivider.clk2[0] ),
    .C(\clkdivider.clk2[2] ),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _0551_ (.A(\clkdivider.clk2[3] ),
    .B(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__nand2_1 _0552_ (.A(\clkdivider.clk2[4] ),
    .B(_0083_),
    .Y(_0084_));
 sky130_fd_sc_hd__or2_1 _0553_ (.A(\clkdivider.clk2[5] ),
    .B(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__xnor2_1 _0554_ (.A(net29),
    .B(_0085_),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _0555_ (.A(\dither.count[0] ),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _0556_ (.A(\stanley.en3[3] ),
    .Y(_0086_));
 sky130_fd_sc_hd__or3_2 _0557_ (.A(\stanley.en3[2] ),
    .B(\stanley.en3[1] ),
    .C(\stanley.en3[0] ),
    .X(_0087_));
 sky130_fd_sc_hd__o21ai_1 _0558_ (.A1(\stanley.en3[1] ),
    .A2(\stanley.en3[0] ),
    .B1(\stanley.en3[2] ),
    .Y(_0088_));
 sky130_fd_sc_hd__and3_1 _0559_ (.A(_0086_),
    .B(_0087_),
    .C(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__clkbuf_2 _0560_ (.A(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__nand2_4 _0561_ (.A(\stanley.en2[3] ),
    .B(\stanley.en2[2] ),
    .Y(_0091_));
 sky130_fd_sc_hd__xnor2_1 _0562_ (.A(\stanley.d_n_1[5] ),
    .B(_0090_),
    .Y(_0092_));
 sky130_fd_sc_hd__nor2_1 _0563_ (.A(_0091_),
    .B(_0092_),
    .Y(_0093_));
 sky130_fd_sc_hd__a21o_1 _0564_ (.A1(\stanley.d_n_1[5] ),
    .A2(_0090_),
    .B1(_0093_),
    .X(_0094_));
 sky130_fd_sc_hd__xor2_1 _0565_ (.A(\stanley.d_n_1[6] ),
    .B(_0090_),
    .X(_0095_));
 sky130_fd_sc_hd__xnor2_1 _0566_ (.A(_0091_),
    .B(_0095_),
    .Y(_0096_));
 sky130_fd_sc_hd__nand2_1 _0567_ (.A(_0094_),
    .B(_0096_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand2_2 _0568_ (.A(net13),
    .B(\stanley.en1[2] ),
    .Y(_0098_));
 sky130_fd_sc_hd__clkbuf_4 _0569_ (.A(_0098_),
    .X(_0099_));
 sky130_fd_sc_hd__xnor2_1 _0570_ (.A(_0094_),
    .B(_0096_),
    .Y(_0100_));
 sky130_fd_sc_hd__or2_1 _0571_ (.A(_0099_),
    .B(_0100_),
    .X(_0101_));
 sky130_fd_sc_hd__and2_1 _0572_ (.A(\stanley.en2[3] ),
    .B(\stanley.en2[2] ),
    .X(_0102_));
 sky130_fd_sc_hd__clkbuf_4 _0573_ (.A(_0102_),
    .X(_0103_));
 sky130_fd_sc_hd__and2_1 _0574_ (.A(\stanley.d_n_1[6] ),
    .B(_0090_),
    .X(_0104_));
 sky130_fd_sc_hd__a21o_1 _0575_ (.A1(_0103_),
    .A2(_0095_),
    .B1(_0104_),
    .X(_0105_));
 sky130_fd_sc_hd__and4_1 _0576_ (.A(_0086_),
    .B(\stanley.d_n_1[7] ),
    .C(_0087_),
    .D(_0088_),
    .X(_0106_));
 sky130_fd_sc_hd__a31o_1 _0577_ (.A1(_0086_),
    .A2(_0087_),
    .A3(_0088_),
    .B1(\stanley.d_n_1[7] ),
    .X(_0107_));
 sky130_fd_sc_hd__or2b_1 _0578_ (.A(_0106_),
    .B_N(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__xnor2_1 _0579_ (.A(_0103_),
    .B(_0108_),
    .Y(_0109_));
 sky130_fd_sc_hd__xnor2_1 _0580_ (.A(_0105_),
    .B(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__or2_1 _0581_ (.A(_0099_),
    .B(_0110_),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_1 _0582_ (.A(_0099_),
    .B(_0110_),
    .Y(_0112_));
 sky130_fd_sc_hd__and2_1 _0583_ (.A(_0111_),
    .B(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__a21bo_1 _0584_ (.A1(_0097_),
    .A2(_0101_),
    .B1_N(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__nand2_1 _0585_ (.A(_0097_),
    .B(_0101_),
    .Y(_0115_));
 sky130_fd_sc_hd__or2_1 _0586_ (.A(_0115_),
    .B(_0113_),
    .X(_0116_));
 sky130_fd_sc_hd__and2_1 _0587_ (.A(_0114_),
    .B(_0116_),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_2 _0588_ (.A(_0117_),
    .X(_0118_));
 sky130_fd_sc_hd__xnor2_1 _0589_ (.A(\stanley.d_n_1[4] ),
    .B(_0090_),
    .Y(_0119_));
 sky130_fd_sc_hd__nand2_1 _0590_ (.A(\stanley.d_n_1[4] ),
    .B(_0090_),
    .Y(_0120_));
 sky130_fd_sc_hd__o21ai_1 _0591_ (.A1(_0091_),
    .A2(_0119_),
    .B1(_0120_),
    .Y(_0121_));
 sky130_fd_sc_hd__and2_1 _0592_ (.A(_0091_),
    .B(_0092_),
    .X(_0122_));
 sky130_fd_sc_hd__nor2_1 _0593_ (.A(_0093_),
    .B(_0122_),
    .Y(_0123_));
 sky130_fd_sc_hd__xnor2_1 _0594_ (.A(_0121_),
    .B(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__nand2_1 _0595_ (.A(_0121_),
    .B(_0123_),
    .Y(_0125_));
 sky130_fd_sc_hd__o21ai_1 _0596_ (.A1(_0099_),
    .A2(_0124_),
    .B1(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__nand2_1 _0597_ (.A(_0099_),
    .B(_0100_),
    .Y(_0127_));
 sky130_fd_sc_hd__and2_1 _0598_ (.A(_0101_),
    .B(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__or2_1 _0599_ (.A(_0126_),
    .B(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__clkbuf_4 _0600_ (.A(\stanley.en3[1] ),
    .X(_0130_));
 sky130_fd_sc_hd__buf_2 _0601_ (.A(\stanley.en3[0] ),
    .X(_0131_));
 sky130_fd_sc_hd__o22ai_1 _0602_ (.A1(\stanley.en3[3] ),
    .A2(\stanley.en3[2] ),
    .B1(_0130_),
    .B2(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__and3_1 _0603_ (.A(\stanley.d_n_1[3] ),
    .B(_0087_),
    .C(_0132_),
    .X(_0133_));
 sky130_fd_sc_hd__a21oi_1 _0604_ (.A1(_0087_),
    .A2(_0132_),
    .B1(\stanley.d_n_1[3] ),
    .Y(_0134_));
 sky130_fd_sc_hd__or3_1 _0605_ (.A(_0091_),
    .B(_0133_),
    .C(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__or2b_1 _0606_ (.A(_0133_),
    .B_N(_0135_),
    .X(_0136_));
 sky130_fd_sc_hd__xnor2_1 _0607_ (.A(_0103_),
    .B(_0119_),
    .Y(_0137_));
 sky130_fd_sc_hd__xnor2_1 _0608_ (.A(_0136_),
    .B(_0137_),
    .Y(_0138_));
 sky130_fd_sc_hd__nand2_1 _0609_ (.A(_0136_),
    .B(_0137_),
    .Y(_0139_));
 sky130_fd_sc_hd__o21ai_1 _0610_ (.A1(_0099_),
    .A2(_0138_),
    .B1(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__xnor2_1 _0611_ (.A(_0099_),
    .B(_0124_),
    .Y(_0141_));
 sky130_fd_sc_hd__xnor2_1 _0612_ (.A(_0140_),
    .B(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__or2b_1 _0613_ (.A(\stanley.en1[0] ),
    .B_N(\stanley.en1[1] ),
    .X(_0143_));
 sky130_fd_sc_hd__or3b_1 _0614_ (.A(\stanley.en1[0] ),
    .B(\stanley.en1[1] ),
    .C_N(\stanley.en1[2] ),
    .X(_0144_));
 sky130_fd_sc_hd__or2_1 _0615_ (.A(\stanley.en1[2] ),
    .B(_0143_),
    .X(_0145_));
 sky130_fd_sc_hd__a21oi_1 _0616_ (.A1(_0144_),
    .A2(_0145_),
    .B1(net13),
    .Y(_0146_));
 sky130_fd_sc_hd__a31o_2 _0617_ (.A1(net13),
    .A2(\stanley.en1[2] ),
    .A3(_0143_),
    .B1(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__or3b_2 _0618_ (.A(\stanley.en2[1] ),
    .B(\stanley.en2[0] ),
    .C_N(\stanley.en2[2] ),
    .X(_0148_));
 sky130_fd_sc_hd__xor2_2 _0619_ (.A(_0130_),
    .B(\stanley.en3[0] ),
    .X(_0149_));
 sky130_fd_sc_hd__xnor2_2 _0620_ (.A(\stanley.en3[3] ),
    .B(\stanley.en3[2] ),
    .Y(_0150_));
 sky130_fd_sc_hd__and3_1 _0621_ (.A(\stanley.d_n_1[2] ),
    .B(_0149_),
    .C(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__a21oi_1 _0622_ (.A1(_0149_),
    .A2(_0150_),
    .B1(\stanley.d_n_1[2] ),
    .Y(_0152_));
 sky130_fd_sc_hd__a211o_1 _0623_ (.A1(_0148_),
    .A2(_0091_),
    .B1(_0151_),
    .C1(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__a21o_1 _0624_ (.A1(_0131_),
    .A2(_0150_),
    .B1(\stanley.d_n_1[1] ),
    .X(_0154_));
 sky130_fd_sc_hd__nor2_1 _0625_ (.A(\stanley.en2[3] ),
    .B(\stanley.en2[2] ),
    .Y(_0155_));
 sky130_fd_sc_hd__o21a_1 _0626_ (.A1(_0155_),
    .A2(_0103_),
    .B1(\stanley.en2[1] ),
    .X(_0156_));
 sky130_fd_sc_hd__and3_1 _0627_ (.A(_0131_),
    .B(\stanley.d_n_1[1] ),
    .C(_0150_),
    .X(_0157_));
 sky130_fd_sc_hd__a21o_1 _0628_ (.A1(_0154_),
    .A2(_0156_),
    .B1(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__nand2_1 _0629_ (.A(_0148_),
    .B(_0091_),
    .Y(_0159_));
 sky130_fd_sc_hd__o21bai_1 _0630_ (.A1(_0151_),
    .A2(_0152_),
    .B1_N(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__and3_1 _0631_ (.A(_0153_),
    .B(_0158_),
    .C(_0160_),
    .X(_0161_));
 sky130_fd_sc_hd__a21o_1 _0632_ (.A1(_0153_),
    .A2(_0160_),
    .B1(_0158_),
    .X(_0162_));
 sky130_fd_sc_hd__and2b_1 _0633_ (.A_N(_0161_),
    .B(_0162_),
    .X(_0163_));
 sky130_fd_sc_hd__xor2_2 _0634_ (.A(_0147_),
    .B(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__a21oi_1 _0635_ (.A1(_0131_),
    .A2(_0150_),
    .B1(\stanley.d_n_1[1] ),
    .Y(_0165_));
 sky130_fd_sc_hd__or3b_1 _0636_ (.A(_0157_),
    .B(_0165_),
    .C_N(_0156_),
    .X(_0166_));
 sky130_fd_sc_hd__o21bai_1 _0637_ (.A1(_0157_),
    .A2(_0165_),
    .B1_N(_0156_),
    .Y(_0167_));
 sky130_fd_sc_hd__inv_2 _0638_ (.A(\stanley.en1[0] ),
    .Y(_0168_));
 sky130_fd_sc_hd__or3b_2 _0639_ (.A(net13),
    .B(\stanley.en1[2] ),
    .C_N(\stanley.en1[0] ),
    .X(_0169_));
 sky130_fd_sc_hd__o21ai_2 _0640_ (.A1(_0168_),
    .A2(_0098_),
    .B1(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__or2_1 _0641_ (.A(_0155_),
    .B(_0103_),
    .X(_0171_));
 sky130_fd_sc_hd__a21o_1 _0642_ (.A1(\stanley.en2[0] ),
    .A2(_0171_),
    .B1(\stanley.d_n_1[0] ),
    .X(_0172_));
 sky130_fd_sc_hd__and3_1 _0643_ (.A(\stanley.en2[0] ),
    .B(\stanley.d_n_1[0] ),
    .C(_0171_),
    .X(_0173_));
 sky130_fd_sc_hd__a21o_1 _0644_ (.A1(_0170_),
    .A2(_0172_),
    .B1(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__xnor2_1 _0645_ (.A(\stanley.en1[0] ),
    .B(\stanley.en1[1] ),
    .Y(_0175_));
 sky130_fd_sc_hd__or2_1 _0646_ (.A(_0098_),
    .B(_0175_),
    .X(_0176_));
 sky130_fd_sc_hd__or3_1 _0647_ (.A(net13),
    .B(\stanley.en1[2] ),
    .C(_0175_),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_1 _0648_ (.A(_0176_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand2_1 _0649_ (.A(_0166_),
    .B(_0167_),
    .Y(_0179_));
 sky130_fd_sc_hd__xnor2_1 _0650_ (.A(_0179_),
    .B(_0174_),
    .Y(_0180_));
 sky130_fd_sc_hd__a32o_2 _0651_ (.A1(_0166_),
    .A2(_0167_),
    .A3(_0174_),
    .B1(_0178_),
    .B2(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__a21o_1 _0652_ (.A1(_0149_),
    .A2(_0150_),
    .B1(\stanley.d_n_1[2] ),
    .X(_0182_));
 sky130_fd_sc_hd__a21o_1 _0653_ (.A1(_0159_),
    .A2(_0182_),
    .B1(_0151_),
    .X(_0183_));
 sky130_fd_sc_hd__o21ai_1 _0654_ (.A1(_0133_),
    .A2(_0134_),
    .B1(_0091_),
    .Y(_0184_));
 sky130_fd_sc_hd__and3_1 _0655_ (.A(_0135_),
    .B(_0183_),
    .C(_0184_),
    .X(_0185_));
 sky130_fd_sc_hd__or2_1 _0656_ (.A(net13),
    .B(_0144_),
    .X(_0186_));
 sky130_fd_sc_hd__a21bo_1 _0657_ (.A1(_0098_),
    .A2(_0169_),
    .B1_N(\stanley.en1[1] ),
    .X(_0187_));
 sky130_fd_sc_hd__nand2_1 _0658_ (.A(_0186_),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _0659_ (.A(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__a21oi_1 _0660_ (.A1(_0135_),
    .A2(_0184_),
    .B1(_0183_),
    .Y(_0190_));
 sky130_fd_sc_hd__nor3_2 _0661_ (.A(_0185_),
    .B(_0189_),
    .C(_0190_),
    .Y(_0191_));
 sky130_fd_sc_hd__o21a_1 _0662_ (.A1(_0185_),
    .A2(_0190_),
    .B1(_0189_),
    .X(_0192_));
 sky130_fd_sc_hd__a21oi_2 _0663_ (.A1(_0147_),
    .A2(_0162_),
    .B1(_0161_),
    .Y(_0193_));
 sky130_fd_sc_hd__o21ai_2 _0664_ (.A1(_0191_),
    .A2(_0192_),
    .B1(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__nor3_1 _0665_ (.A(_0191_),
    .B(_0193_),
    .C(_0192_),
    .Y(_0195_));
 sky130_fd_sc_hd__a31o_1 _0666_ (.A1(_0164_),
    .A2(_0181_),
    .A3(_0194_),
    .B1(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__nor2_1 _0667_ (.A(_0185_),
    .B(_0191_),
    .Y(_0197_));
 sky130_fd_sc_hd__xor2_1 _0668_ (.A(_0099_),
    .B(_0138_),
    .X(_0198_));
 sky130_fd_sc_hd__xnor2_1 _0669_ (.A(_0197_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__and2b_1 _0670_ (.A_N(_0197_),
    .B(_0198_),
    .X(_0200_));
 sky130_fd_sc_hd__a21o_1 _0671_ (.A1(_0196_),
    .A2(_0199_),
    .B1(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__and2b_1 _0672_ (.A_N(_0141_),
    .B(_0140_),
    .X(_0202_));
 sky130_fd_sc_hd__a21o_1 _0673_ (.A1(_0142_),
    .A2(_0201_),
    .B1(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__and3_1 _0674_ (.A(_0101_),
    .B(_0126_),
    .C(_0127_),
    .X(_0204_));
 sky130_fd_sc_hd__a21o_2 _0675_ (.A1(_0129_),
    .A2(_0203_),
    .B1(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__xor2_2 _0676_ (.A(_0118_),
    .B(_0205_),
    .X(_0206_));
 sky130_fd_sc_hd__nand2_2 _0677_ (.A(\stanley.en[3] ),
    .B(\stanley.en[2] ),
    .Y(_0207_));
 sky130_fd_sc_hd__o21bai_1 _0678_ (.A1(\stanley.en1[0] ),
    .A2(\stanley.en1[1] ),
    .B1_N(\stanley.en1[2] ),
    .Y(_0208_));
 sky130_fd_sc_hd__a21o_2 _0679_ (.A1(_0208_),
    .A2(_0144_),
    .B1(net13),
    .X(_0209_));
 sky130_fd_sc_hd__o21bai_1 _0680_ (.A1(\stanley.en2[1] ),
    .A2(\stanley.en2[0] ),
    .B1_N(\stanley.en2[2] ),
    .Y(_0210_));
 sky130_fd_sc_hd__a21o_2 _0681_ (.A1(_0210_),
    .A2(_0148_),
    .B1(\stanley.en2[3] ),
    .X(_0211_));
 sky130_fd_sc_hd__buf_2 _0682_ (.A(\stanley.en3[3] ),
    .X(_0212_));
 sky130_fd_sc_hd__buf_2 _0683_ (.A(\stanley.en3[2] ),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _0684_ (.A(_0212_),
    .B(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__nand2_1 _0685_ (.A(\stanley.d_n_1[13] ),
    .B(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__or2_1 _0686_ (.A(\stanley.d_n_1[13] ),
    .B(_0214_),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_1 _0687_ (.A(_0215_),
    .B(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__xor2_1 _0688_ (.A(_0211_),
    .B(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__nand2_1 _0689_ (.A(_0212_),
    .B(_0213_),
    .Y(_0219_));
 sky130_fd_sc_hd__nor2_1 _0690_ (.A(_0130_),
    .B(_0131_),
    .Y(_0220_));
 sky130_fd_sc_hd__or4b_1 _0691_ (.A(_0212_),
    .B(_0130_),
    .C(_0131_),
    .D_N(_0213_),
    .X(_0221_));
 sky130_fd_sc_hd__o21ai_2 _0692_ (.A1(_0219_),
    .A2(_0220_),
    .B1(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__xnor2_1 _0693_ (.A(\stanley.d_n_1[12] ),
    .B(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__inv_2 _0694_ (.A(_0155_),
    .Y(_0224_));
 sky130_fd_sc_hd__xnor2_1 _0695_ (.A(\stanley.en2[1] ),
    .B(\stanley.en2[0] ),
    .Y(_0225_));
 sky130_fd_sc_hd__o22a_1 _0696_ (.A1(_0224_),
    .A2(_0225_),
    .B1(_0091_),
    .B2(\stanley.en2[1] ),
    .X(_0226_));
 sky130_fd_sc_hd__nor2_1 _0697_ (.A(_0223_),
    .B(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__a21oi_1 _0698_ (.A1(\stanley.d_n_1[12] ),
    .A2(_0222_),
    .B1(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__xnor2_1 _0699_ (.A(_0218_),
    .B(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__xnor2_1 _0700_ (.A(_0209_),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__and2_1 _0701_ (.A(_0223_),
    .B(_0226_),
    .X(_0231_));
 sky130_fd_sc_hd__or2_1 _0702_ (.A(_0227_),
    .B(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__or3b_1 _0703_ (.A(_0212_),
    .B(_0213_),
    .C_N(_0130_),
    .X(_0233_));
 sky130_fd_sc_hd__o21ai_2 _0704_ (.A1(_0219_),
    .A2(_0149_),
    .B1(_0233_),
    .Y(_0234_));
 sky130_fd_sc_hd__xor2_2 _0705_ (.A(\stanley.d_n_1[11] ),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__inv_2 _0706_ (.A(\stanley.en2[0] ),
    .Y(_0236_));
 sky130_fd_sc_hd__or2b_1 _0707_ (.A(\stanley.en2[2] ),
    .B_N(\stanley.en2[0] ),
    .X(_0237_));
 sky130_fd_sc_hd__a21oi_1 _0708_ (.A1(_0148_),
    .A2(_0237_),
    .B1(\stanley.en2[3] ),
    .Y(_0238_));
 sky130_fd_sc_hd__a31o_1 _0709_ (.A1(\stanley.en2[1] ),
    .A2(_0236_),
    .A3(_0103_),
    .B1(_0238_),
    .X(_0239_));
 sky130_fd_sc_hd__and2_1 _0710_ (.A(\stanley.d_n_1[11] ),
    .B(_0234_),
    .X(_0240_));
 sky130_fd_sc_hd__a21o_1 _0711_ (.A1(_0235_),
    .A2(_0239_),
    .B1(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__xor2_1 _0712_ (.A(_0232_),
    .B(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__o32a_1 _0713_ (.A1(\stanley.en1[0] ),
    .A2(\stanley.en1[1] ),
    .A3(_0099_),
    .B1(_0208_),
    .B2(net13),
    .X(_0243_));
 sky130_fd_sc_hd__or2b_1 _0714_ (.A(_0232_),
    .B_N(_0241_),
    .X(_0244_));
 sky130_fd_sc_hd__o21a_1 _0715_ (.A1(_0242_),
    .A2(_0243_),
    .B1(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__xor2_1 _0716_ (.A(_0230_),
    .B(_0245_),
    .X(_0246_));
 sky130_fd_sc_hd__nor2_1 _0717_ (.A(_0207_),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__and2_1 _0718_ (.A(_0207_),
    .B(_0246_),
    .X(_0248_));
 sky130_fd_sc_hd__nor2_1 _0719_ (.A(_0247_),
    .B(_0248_),
    .Y(_0249_));
 sky130_fd_sc_hd__xnor2_1 _0720_ (.A(_0242_),
    .B(_0243_),
    .Y(_0250_));
 sky130_fd_sc_hd__or4_1 _0721_ (.A(\stanley.en1[3] ),
    .B(\stanley.en1[2] ),
    .C(_0168_),
    .D(\stanley.en1[1] ),
    .X(_0251_));
 sky130_fd_sc_hd__and3_1 _0722_ (.A(_0186_),
    .B(_0176_),
    .C(_0251_),
    .X(_0252_));
 sky130_fd_sc_hd__or3b_1 _0723_ (.A(_0212_),
    .B(\stanley.en3[2] ),
    .C_N(_0131_),
    .X(_0253_));
 sky130_fd_sc_hd__nand3b_1 _0724_ (.A_N(_0131_),
    .B(_0213_),
    .C(_0212_),
    .Y(_0254_));
 sky130_fd_sc_hd__inv_2 _0725_ (.A(\stanley.d_n_1[10] ),
    .Y(_0255_));
 sky130_fd_sc_hd__a21o_1 _0726_ (.A1(_0253_),
    .A2(_0254_),
    .B1(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__a22o_1 _0727_ (.A1(\stanley.en2[1] ),
    .A2(_0155_),
    .B1(_0225_),
    .B2(_0103_),
    .X(_0257_));
 sky130_fd_sc_hd__nand3_1 _0728_ (.A(_0255_),
    .B(_0253_),
    .C(_0254_),
    .Y(_0258_));
 sky130_fd_sc_hd__nand3_1 _0729_ (.A(_0256_),
    .B(_0257_),
    .C(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__nand2_1 _0730_ (.A(_0256_),
    .B(_0259_),
    .Y(_0260_));
 sky130_fd_sc_hd__xor2_2 _0731_ (.A(_0235_),
    .B(_0239_),
    .X(_0261_));
 sky130_fd_sc_hd__xnor2_2 _0732_ (.A(_0260_),
    .B(_0261_),
    .Y(_0262_));
 sky130_fd_sc_hd__nand2_1 _0733_ (.A(_0260_),
    .B(_0261_),
    .Y(_0263_));
 sky130_fd_sc_hd__o21ai_1 _0734_ (.A1(_0252_),
    .A2(_0262_),
    .B1(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__and2b_1 _0735_ (.A_N(_0250_),
    .B(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__inv_2 _0736_ (.A(\stanley.en[3] ),
    .Y(_0266_));
 sky130_fd_sc_hd__or2_1 _0737_ (.A(\stanley.en[0] ),
    .B(\stanley.en[1] ),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_1 _0738_ (.A(\stanley.en[2] ),
    .B(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__a21o_1 _0739_ (.A1(\stanley.en[0] ),
    .A2(\stanley.en[1] ),
    .B1(\stanley.en[2] ),
    .X(_0269_));
 sky130_fd_sc_hd__and2_1 _0740_ (.A(\stanley.en[3] ),
    .B(\stanley.en[2] ),
    .X(_0270_));
 sky130_fd_sc_hd__buf_2 _0741_ (.A(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__a32o_1 _0742_ (.A1(_0266_),
    .A2(_0268_),
    .A3(_0269_),
    .B1(\stanley.en[1] ),
    .B2(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__xnor2_1 _0743_ (.A(_0264_),
    .B(_0250_),
    .Y(_0273_));
 sky130_fd_sc_hd__and2_1 _0744_ (.A(_0272_),
    .B(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__nor3_1 _0745_ (.A(_0249_),
    .B(_0265_),
    .C(_0274_),
    .Y(_0275_));
 sky130_fd_sc_hd__o21a_1 _0746_ (.A1(_0265_),
    .A2(_0274_),
    .B1(_0249_),
    .X(_0276_));
 sky130_fd_sc_hd__or2_1 _0747_ (.A(_0275_),
    .B(_0276_),
    .X(_0277_));
 sky130_fd_sc_hd__xnor2_1 _0748_ (.A(_0272_),
    .B(_0273_),
    .Y(_0278_));
 sky130_fd_sc_hd__a21bo_1 _0749_ (.A1(_0213_),
    .A2(_0130_),
    .B1_N(_0212_),
    .X(_0279_));
 sky130_fd_sc_hd__nand3b_2 _0750_ (.A_N(\stanley.en3[3] ),
    .B(_0213_),
    .C(_0130_),
    .Y(_0280_));
 sky130_fd_sc_hd__mux2_1 _0751_ (.A0(_0213_),
    .A1(_0130_),
    .S(\stanley.en3[0] ),
    .X(_0281_));
 sky130_fd_sc_hd__a31o_1 _0752_ (.A1(_0279_),
    .A2(_0280_),
    .A3(_0281_),
    .B1(\stanley.d_n_1[9] ),
    .X(_0282_));
 sky130_fd_sc_hd__a2bb2o_1 _0753_ (.A1_N(\stanley.en2[3] ),
    .A2_N(_0237_),
    .B1(_0236_),
    .B2(_0102_),
    .X(_0283_));
 sky130_fd_sc_hd__nand4_1 _0754_ (.A(\stanley.d_n_1[9] ),
    .B(_0279_),
    .C(_0280_),
    .D(_0281_),
    .Y(_0284_));
 sky130_fd_sc_hd__a21bo_1 _0755_ (.A1(_0282_),
    .A2(_0283_),
    .B1_N(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__a21o_1 _0756_ (.A1(_0256_),
    .A2(_0258_),
    .B1(_0257_),
    .X(_0286_));
 sky130_fd_sc_hd__nand3_1 _0757_ (.A(_0259_),
    .B(_0285_),
    .C(_0286_),
    .Y(_0287_));
 sky130_fd_sc_hd__a31o_1 _0758_ (.A1(net13),
    .A2(\stanley.en1[2] ),
    .A3(\stanley.en1[0] ),
    .B1(_0146_),
    .X(_0288_));
 sky130_fd_sc_hd__a21o_1 _0759_ (.A1(_0259_),
    .A2(_0286_),
    .B1(_0285_),
    .X(_0289_));
 sky130_fd_sc_hd__and3_1 _0760_ (.A(_0287_),
    .B(_0288_),
    .C(_0289_),
    .X(_0290_));
 sky130_fd_sc_hd__a31o_1 _0761_ (.A1(_0259_),
    .A2(_0285_),
    .A3(_0286_),
    .B1(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__xor2_2 _0762_ (.A(_0252_),
    .B(_0262_),
    .X(_0292_));
 sky130_fd_sc_hd__xnor2_2 _0763_ (.A(_0291_),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _0764_ (.A(\stanley.en[0] ),
    .Y(_0294_));
 sky130_fd_sc_hd__nor2_1 _0765_ (.A(\stanley.en[3] ),
    .B(\stanley.en[2] ),
    .Y(_0295_));
 sky130_fd_sc_hd__o21ai_1 _0766_ (.A1(_0266_),
    .A2(_0294_),
    .B1(_0267_),
    .Y(_0296_));
 sky130_fd_sc_hd__a32o_1 _0767_ (.A1(_0294_),
    .A2(\stanley.en[1] ),
    .A3(_0295_),
    .B1(_0296_),
    .B2(\stanley.en[2] ),
    .X(_0297_));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__o2bb2a_1 _0769_ (.A1_N(_0291_),
    .A2_N(_0292_),
    .B1(_0293_),
    .B2(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__or2_1 _0770_ (.A(_0278_),
    .B(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__xnor2_2 _0771_ (.A(_0293_),
    .B(_0297_),
    .Y(_0301_));
 sky130_fd_sc_hd__o21ai_2 _0772_ (.A1(\stanley.en1[1] ),
    .A2(_0098_),
    .B1(_0177_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand3_1 _0773_ (.A(_0284_),
    .B(_0282_),
    .C(_0283_),
    .Y(_0303_));
 sky130_fd_sc_hd__a21o_1 _0774_ (.A1(_0284_),
    .A2(_0282_),
    .B1(_0283_),
    .X(_0304_));
 sky130_fd_sc_hd__a21bo_1 _0775_ (.A1(\stanley.en3[2] ),
    .A2(_0131_),
    .B1_N(\stanley.en3[3] ),
    .X(_0305_));
 sky130_fd_sc_hd__or2_1 _0776_ (.A(\stanley.en3[2] ),
    .B(_0130_),
    .X(_0306_));
 sky130_fd_sc_hd__or2b_1 _0777_ (.A(\stanley.en3[3] ),
    .B_N(_0131_),
    .X(_0307_));
 sky130_fd_sc_hd__a41o_1 _0778_ (.A1(_0280_),
    .A2(_0305_),
    .A3(_0306_),
    .A4(_0307_),
    .B1(\stanley.d_n_1[8] ),
    .X(_0308_));
 sky130_fd_sc_hd__o21ba_1 _0779_ (.A1(_0213_),
    .A2(_0130_),
    .B1_N(\stanley.en3[0] ),
    .X(_0309_));
 sky130_fd_sc_hd__o2111a_1 _0780_ (.A1(_0212_),
    .A2(_0309_),
    .B1(_0305_),
    .C1(_0280_),
    .D1(\stanley.d_n_1[8] ),
    .X(_0310_));
 sky130_fd_sc_hd__a21o_1 _0781_ (.A1(_0103_),
    .A2(_0308_),
    .B1(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__a21o_1 _0782_ (.A1(_0303_),
    .A2(_0304_),
    .B1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__nand3_1 _0783_ (.A(_0303_),
    .B(_0311_),
    .C(_0304_),
    .Y(_0313_));
 sky130_fd_sc_hd__a21boi_2 _0784_ (.A1(_0302_),
    .A2(_0312_),
    .B1_N(_0313_),
    .Y(_0314_));
 sky130_fd_sc_hd__a21oi_1 _0785_ (.A1(_0287_),
    .A2(_0289_),
    .B1(_0288_),
    .Y(_0315_));
 sky130_fd_sc_hd__nor2_1 _0786_ (.A(_0290_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__xnor2_2 _0787_ (.A(_0314_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand2_1 _0788_ (.A(\stanley.en[0] ),
    .B(\stanley.en[1] ),
    .Y(_0318_));
 sky130_fd_sc_hd__o211a_1 _0789_ (.A1(_0271_),
    .A2(_0295_),
    .B1(_0318_),
    .C1(_0267_),
    .X(_0319_));
 sky130_fd_sc_hd__or3_1 _0790_ (.A(_0290_),
    .B(_0314_),
    .C(_0315_),
    .X(_0320_));
 sky130_fd_sc_hd__a21boi_2 _0791_ (.A1(_0317_),
    .A2(_0319_),
    .B1_N(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__xnor2_2 _0792_ (.A(_0301_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__xnor2_2 _0793_ (.A(_0317_),
    .B(_0319_),
    .Y(_0323_));
 sky130_fd_sc_hd__o21ai_2 _0794_ (.A1(_0271_),
    .A2(_0295_),
    .B1(\stanley.en[0] ),
    .Y(_0324_));
 sky130_fd_sc_hd__and3_1 _0795_ (.A(_0313_),
    .B(_0302_),
    .C(_0312_),
    .X(_0325_));
 sky130_fd_sc_hd__o21ai_2 _0796_ (.A1(\stanley.en1[0] ),
    .A2(_0099_),
    .B1(_0169_),
    .Y(_0326_));
 sky130_fd_sc_hd__or3b_1 _0797_ (.A(_0091_),
    .B(_0310_),
    .C_N(_0308_),
    .X(_0327_));
 sky130_fd_sc_hd__o2111ai_1 _0798_ (.A1(_0212_),
    .A2(_0309_),
    .B1(_0305_),
    .C1(_0280_),
    .D1(\stanley.d_n_1[8] ),
    .Y(_0328_));
 sky130_fd_sc_hd__a21o_1 _0799_ (.A1(_0328_),
    .A2(_0308_),
    .B1(_0103_),
    .X(_0329_));
 sky130_fd_sc_hd__a21o_1 _0800_ (.A1(_0103_),
    .A2(_0107_),
    .B1(_0106_),
    .X(_0330_));
 sky130_fd_sc_hd__a21o_1 _0801_ (.A1(_0327_),
    .A2(_0329_),
    .B1(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__and3_1 _0802_ (.A(_0327_),
    .B(_0330_),
    .C(_0329_),
    .X(_0332_));
 sky130_fd_sc_hd__a21oi_1 _0803_ (.A1(_0326_),
    .A2(_0331_),
    .B1(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__a21oi_1 _0804_ (.A1(_0313_),
    .A2(_0312_),
    .B1(_0302_),
    .Y(_0334_));
 sky130_fd_sc_hd__or3_1 _0805_ (.A(_0325_),
    .B(_0333_),
    .C(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__o21ai_1 _0806_ (.A1(_0325_),
    .A2(_0334_),
    .B1(_0333_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand2_1 _0807_ (.A(_0335_),
    .B(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__o21ai_2 _0808_ (.A1(_0324_),
    .A2(_0337_),
    .B1(_0335_),
    .Y(_0338_));
 sky130_fd_sc_hd__xnor2_2 _0809_ (.A(_0323_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__and2_1 _0810_ (.A(_0322_),
    .B(_0339_),
    .X(_0340_));
 sky130_fd_sc_hd__nand2_1 _0811_ (.A(_0105_),
    .B(_0109_),
    .Y(_0341_));
 sky130_fd_sc_hd__and2b_1 _0812_ (.A_N(_0332_),
    .B(_0331_),
    .X(_0342_));
 sky130_fd_sc_hd__xnor2_1 _0813_ (.A(_0326_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__a21oi_1 _0814_ (.A1(_0341_),
    .A2(_0111_),
    .B1(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__and3_1 _0815_ (.A(_0341_),
    .B(_0111_),
    .C(_0343_),
    .X(_0345_));
 sky130_fd_sc_hd__or2_1 _0816_ (.A(_0344_),
    .B(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__nor2_1 _0817_ (.A(_0114_),
    .B(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__xor2_1 _0818_ (.A(_0324_),
    .B(_0337_),
    .X(_0348_));
 sky130_fd_sc_hd__o21a_1 _0819_ (.A1(_0344_),
    .A2(_0347_),
    .B1(_0348_),
    .X(_0349_));
 sky130_fd_sc_hd__and2_1 _0820_ (.A(_0340_),
    .B(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__xnor2_1 _0821_ (.A(_0348_),
    .B(_0344_),
    .Y(_0351_));
 sky130_fd_sc_hd__xor2_1 _0822_ (.A(_0114_),
    .B(_0346_),
    .X(_0352_));
 sky130_fd_sc_hd__and2b_1 _0823_ (.A_N(_0351_),
    .B(_0352_),
    .X(_0353_));
 sky130_fd_sc_hd__and4_1 _0824_ (.A(_0340_),
    .B(_0118_),
    .C(_0205_),
    .D(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__or2b_1 _0825_ (.A(_0301_),
    .B_N(_0321_),
    .X(_0355_));
 sky130_fd_sc_hd__and2b_1 _0826_ (.A_N(_0323_),
    .B(_0338_),
    .X(_0356_));
 sky130_fd_sc_hd__and2b_1 _0827_ (.A_N(_0321_),
    .B(_0301_),
    .X(_0357_));
 sky130_fd_sc_hd__a21o_1 _0828_ (.A1(_0355_),
    .A2(_0356_),
    .B1(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__nand2_1 _0829_ (.A(_0278_),
    .B(_0299_),
    .Y(_0359_));
 sky130_fd_sc_hd__and2_1 _0830_ (.A(_0300_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__o31ai_4 _0831_ (.A1(_0350_),
    .A2(_0354_),
    .A3(_0358_),
    .B1(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2_1 _0832_ (.A(_0300_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__xnor2_2 _0833_ (.A(_0277_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__nand2_1 _0834_ (.A(\stanley.d_n_1[14] ),
    .B(_0214_),
    .Y(_0364_));
 sky130_fd_sc_hd__nor2_1 _0835_ (.A(\stanley.d_n_1[14] ),
    .B(_0214_),
    .Y(_0365_));
 sky130_fd_sc_hd__inv_2 _0836_ (.A(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__nand2_1 _0837_ (.A(_0364_),
    .B(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__xnor2_1 _0838_ (.A(_0211_),
    .B(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__o21ai_1 _0839_ (.A1(_0211_),
    .A2(_0217_),
    .B1(_0215_),
    .Y(_0369_));
 sky130_fd_sc_hd__xnor2_1 _0840_ (.A(_0368_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__and2b_1 _0841_ (.A_N(_0209_),
    .B(_0370_),
    .X(_0371_));
 sky130_fd_sc_hd__and2b_1 _0842_ (.A_N(_0370_),
    .B(_0209_),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _0843_ (.A(_0371_),
    .B(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__inv_2 _0844_ (.A(_0229_),
    .Y(_0374_));
 sky130_fd_sc_hd__or2b_1 _0845_ (.A(_0228_),
    .B_N(_0218_),
    .X(_0375_));
 sky130_fd_sc_hd__o21a_1 _0846_ (.A1(_0209_),
    .A2(_0374_),
    .B1(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__xnor2_1 _0847_ (.A(_0373_),
    .B(_0376_),
    .Y(_0377_));
 sky130_fd_sc_hd__xnor2_1 _0848_ (.A(_0271_),
    .B(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__and2b_1 _0849_ (.A_N(_0245_),
    .B(_0230_),
    .X(_0379_));
 sky130_fd_sc_hd__nor2_1 _0850_ (.A(_0379_),
    .B(_0247_),
    .Y(_0380_));
 sky130_fd_sc_hd__xnor2_1 _0851_ (.A(_0378_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__inv_2 _0852_ (.A(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__o21ba_1 _0853_ (.A1(_0278_),
    .A2(_0299_),
    .B1_N(_0276_),
    .X(_0383_));
 sky130_fd_sc_hd__a21oi_1 _0854_ (.A1(_0383_),
    .A2(_0361_),
    .B1(_0275_),
    .Y(_0384_));
 sky130_fd_sc_hd__xnor2_2 _0855_ (.A(_0382_),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__a31o_1 _0856_ (.A1(_0118_),
    .A2(_0205_),
    .A3(_0353_),
    .B1(_0349_),
    .X(_0386_));
 sky130_fd_sc_hd__a21o_1 _0857_ (.A1(_0339_),
    .A2(_0386_),
    .B1(_0356_),
    .X(_0387_));
 sky130_fd_sc_hd__xnor2_2 _0858_ (.A(_0322_),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__xnor2_1 _0859_ (.A(_0339_),
    .B(_0386_),
    .Y(_0389_));
 sky130_fd_sc_hd__or3_1 _0860_ (.A(_0191_),
    .B(_0193_),
    .C(_0192_),
    .X(_0390_));
 sky130_fd_sc_hd__and4_1 _0861_ (.A(_0390_),
    .B(_0164_),
    .C(_0181_),
    .D(_0194_),
    .X(_0391_));
 sky130_fd_sc_hd__a22oi_2 _0862_ (.A1(_0164_),
    .A2(_0181_),
    .B1(_0194_),
    .B2(_0390_),
    .Y(_0392_));
 sky130_fd_sc_hd__xnor2_1 _0863_ (.A(_0164_),
    .B(_0181_),
    .Y(_0393_));
 sky130_fd_sc_hd__xnor2_1 _0864_ (.A(_0178_),
    .B(_0180_),
    .Y(_0394_));
 sky130_fd_sc_hd__or2_1 _0865_ (.A(_0393_),
    .B(_0394_),
    .X(_0395_));
 sky130_fd_sc_hd__xnor2_1 _0866_ (.A(_0142_),
    .B(_0201_),
    .Y(_0396_));
 sky130_fd_sc_hd__xnor2_1 _0867_ (.A(_0196_),
    .B(_0199_),
    .Y(_0397_));
 sky130_fd_sc_hd__o311a_1 _0868_ (.A1(_0391_),
    .A2(_0392_),
    .A3(_0395_),
    .B1(_0396_),
    .C1(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__and2b_1 _0869_ (.A_N(_0204_),
    .B(_0129_),
    .X(_0399_));
 sky130_fd_sc_hd__xnor2_2 _0870_ (.A(_0399_),
    .B(_0203_),
    .Y(_0400_));
 sky130_fd_sc_hd__or3b_1 _0871_ (.A(_0398_),
    .B(_0400_),
    .C_N(_0206_),
    .X(_0401_));
 sky130_fd_sc_hd__inv_2 _0872_ (.A(_0346_),
    .Y(_0402_));
 sky130_fd_sc_hd__a21oi_1 _0873_ (.A1(_0118_),
    .A2(_0205_),
    .B1(_0352_),
    .Y(_0403_));
 sky130_fd_sc_hd__a31o_1 _0874_ (.A1(_0402_),
    .A2(_0118_),
    .A3(_0205_),
    .B1(_0403_),
    .X(_0404_));
 sky130_fd_sc_hd__a31o_1 _0875_ (.A1(_0402_),
    .A2(_0118_),
    .A3(_0205_),
    .B1(_0347_),
    .X(_0405_));
 sky130_fd_sc_hd__xor2_1 _0876_ (.A(_0351_),
    .B(_0405_),
    .X(_0406_));
 sky130_fd_sc_hd__nand4_1 _0877_ (.A(_0389_),
    .B(_0401_),
    .C(_0404_),
    .D(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__or4_1 _0878_ (.A(_0350_),
    .B(_0354_),
    .C(_0358_),
    .D(_0360_),
    .X(_0408_));
 sky130_fd_sc_hd__and4b_1 _0879_ (.A_N(_0388_),
    .B(_0407_),
    .C(_0408_),
    .D(_0361_),
    .X(_0409_));
 sky130_fd_sc_hd__and3_2 _0880_ (.A(_0363_),
    .B(_0385_),
    .C(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__or2b_1 _0881_ (.A(_0380_),
    .B_N(_0378_),
    .X(_0411_));
 sky130_fd_sc_hd__a211o_1 _0882_ (.A1(_0383_),
    .A2(_0361_),
    .B1(_0382_),
    .C1(_0275_),
    .X(_0412_));
 sky130_fd_sc_hd__and2b_1 _0883_ (.A_N(_0368_),
    .B(_0369_),
    .X(_0413_));
 sky130_fd_sc_hd__o21a_1 _0884_ (.A1(_0211_),
    .A2(_0365_),
    .B1(_0364_),
    .X(_0414_));
 sky130_fd_sc_hd__nor2_1 _0885_ (.A(\stanley.d_n_1[15] ),
    .B(_0214_),
    .Y(_0415_));
 sky130_fd_sc_hd__and3_1 _0886_ (.A(_0212_),
    .B(_0213_),
    .C(\stanley.d_n_1[15] ),
    .X(_0416_));
 sky130_fd_sc_hd__or2_1 _0887_ (.A(_0415_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__xnor2_1 _0888_ (.A(_0211_),
    .B(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__nor2_1 _0889_ (.A(_0414_),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__and2_1 _0890_ (.A(_0414_),
    .B(_0418_),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_1 _0891_ (.A(_0419_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__xnor2_1 _0892_ (.A(_0421_),
    .B(_0209_),
    .Y(_0422_));
 sky130_fd_sc_hd__o21a_1 _0893_ (.A1(_0413_),
    .A2(_0371_),
    .B1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__nor3_1 _0894_ (.A(_0422_),
    .B(_0413_),
    .C(_0371_),
    .Y(_0424_));
 sky130_fd_sc_hd__nor2_1 _0895_ (.A(_0423_),
    .B(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__xnor2_1 _0896_ (.A(_0207_),
    .B(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__nor2_1 _0897_ (.A(_0373_),
    .B(_0376_),
    .Y(_0427_));
 sky130_fd_sc_hd__nor2_1 _0898_ (.A(_0207_),
    .B(_0377_),
    .Y(_0428_));
 sky130_fd_sc_hd__nor3_1 _0899_ (.A(_0426_),
    .B(_0427_),
    .C(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__o21a_1 _0900_ (.A1(_0427_),
    .A2(_0428_),
    .B1(_0426_),
    .X(_0430_));
 sky130_fd_sc_hd__or2_1 _0901_ (.A(_0429_),
    .B(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__nand3_2 _0902_ (.A(_0411_),
    .B(_0412_),
    .C(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__a21o_1 _0903_ (.A1(_0411_),
    .A2(_0412_),
    .B1(_0431_),
    .X(_0433_));
 sky130_fd_sc_hd__and2_1 _0904_ (.A(_0432_),
    .B(_0433_),
    .X(_0434_));
 sky130_fd_sc_hd__buf_2 _0905_ (.A(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__a21o_1 _0906_ (.A1(_0271_),
    .A2(_0425_),
    .B1(_0423_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_1 _0907_ (.A0(_0416_),
    .A1(_0415_),
    .S(_0211_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _0908_ (.A0(_0420_),
    .A1(_0419_),
    .S(_0209_),
    .X(_0438_));
 sky130_fd_sc_hd__xor2_2 _0909_ (.A(_0437_),
    .B(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__xnor2_2 _0910_ (.A(_0271_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__xnor2_4 _0911_ (.A(_0436_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__inv_2 _0912_ (.A(_0430_),
    .Y(_0442_));
 sky130_fd_sc_hd__a31o_2 _0913_ (.A1(_0442_),
    .A2(_0411_),
    .A3(_0412_),
    .B1(_0429_),
    .X(_0443_));
 sky130_fd_sc_hd__xnor2_4 _0914_ (.A(_0441_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__o31a_1 _0915_ (.A1(_0206_),
    .A2(_0410_),
    .A3(_0435_),
    .B1(_0444_),
    .X(\dither.d_n_input[1] ));
 sky130_fd_sc_hd__xor2_4 _0916_ (.A(_0441_),
    .B(_0443_),
    .X(_0445_));
 sky130_fd_sc_hd__o41ai_1 _0917_ (.A1(_0445_),
    .A2(_0404_),
    .A3(_0410_),
    .A4(_0435_),
    .B1(_0008_),
    .Y(_0446_));
 sky130_fd_sc_hd__o311a_1 _0918_ (.A1(\dither.count[1] ),
    .A2(_0008_),
    .A3(\dither.d_n_input[1] ),
    .B1(_0446_),
    .C1(\dither.count[2] ),
    .X(_0447_));
 sky130_fd_sc_hd__o311ai_4 _0919_ (.A1(_0206_),
    .A2(_0410_),
    .A3(_0435_),
    .B1(_0444_),
    .C1(\dither.count[1] ),
    .Y(_0448_));
 sky130_fd_sc_hd__nor3_1 _0920_ (.A(\dither.count[0] ),
    .B(\dither.count[2] ),
    .C(_0448_),
    .Y(_0449_));
 sky130_fd_sc_hd__a32oi_4 _0921_ (.A1(_0363_),
    .A2(_0385_),
    .A3(_0409_),
    .B1(_0432_),
    .B2(_0433_),
    .Y(_0450_));
 sky130_fd_sc_hd__a21oi_2 _0922_ (.A1(_0400_),
    .A2(_0450_),
    .B1(_0445_),
    .Y(\dither.d_n_input[0] ));
 sky130_fd_sc_hd__o21ai_2 _0923_ (.A1(_0447_),
    .A2(_0449_),
    .B1(\dither.d_n_input[0] ),
    .Y(_0451_));
 sky130_fd_sc_hd__inv_2 _0924_ (.A(_0400_),
    .Y(_0452_));
 sky130_fd_sc_hd__nand2_4 _0925_ (.A(_0444_),
    .B(_0450_),
    .Y(_0453_));
 sky130_fd_sc_hd__o311a_1 _0926_ (.A1(_0452_),
    .A2(_0410_),
    .A3(_0435_),
    .B1(_0444_),
    .C1(\dither.count[2] ),
    .X(_0454_));
 sky130_fd_sc_hd__or3b_2 _0927_ (.A(_0445_),
    .B(_0404_),
    .C_N(_0450_),
    .X(_0455_));
 sky130_fd_sc_hd__o32ai_4 _0928_ (.A1(_0452_),
    .A2(_0453_),
    .A3(_0448_),
    .B1(_0454_),
    .B2(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__nor2_1 _0929_ (.A(_0455_),
    .B(_0448_),
    .Y(_0457_));
 sky130_fd_sc_hd__a21oi_2 _0930_ (.A1(\dither.count[0] ),
    .A2(_0456_),
    .B1(_0457_),
    .Y(_0458_));
 sky130_fd_sc_hd__or2_2 _0931_ (.A(_0406_),
    .B(_0453_),
    .X(_0459_));
 sky130_fd_sc_hd__a21oi_2 _0932_ (.A1(_0451_),
    .A2(_0458_),
    .B1(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__nor2_1 _0933_ (.A(_0389_),
    .B(_0453_),
    .Y(\dither.d_n_input[4] ));
 sky130_fd_sc_hd__a21oi_4 _0934_ (.A1(_0388_),
    .A2(_0450_),
    .B1(_0445_),
    .Y(\dither.d_n_input[5] ));
 sky130_fd_sc_hd__a211o_2 _0935_ (.A1(_0451_),
    .A2(_0458_),
    .B1(_0459_),
    .C1(_0389_),
    .X(_0461_));
 sky130_fd_sc_hd__o211ai_4 _0936_ (.A1(_0460_),
    .A2(\dither.d_n_input[4] ),
    .B1(\dither.d_n_input[5] ),
    .C1(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__a21o_1 _0937_ (.A1(_0361_),
    .A2(_0408_),
    .B1(_0453_),
    .X(_0463_));
 sky130_fd_sc_hd__and2_1 _0938_ (.A(_0444_),
    .B(_0463_),
    .X(_0464_));
 sky130_fd_sc_hd__buf_1 _0939_ (.A(_0464_),
    .X(\dither.d_n_input[6] ));
 sky130_fd_sc_hd__inv_2 _0940_ (.A(\dither.d_n_input[6] ),
    .Y(_0465_));
 sky130_fd_sc_hd__o21a_1 _0941_ (.A1(_0447_),
    .A2(_0449_),
    .B1(\dither.d_n_input[0] ),
    .X(_0466_));
 sky130_fd_sc_hd__a21o_1 _0942_ (.A1(\dither.count[0] ),
    .A2(_0456_),
    .B1(_0457_),
    .X(_0467_));
 sky130_fd_sc_hd__inv_2 _0943_ (.A(_0459_),
    .Y(\dither.d_n_input[3] ));
 sky130_fd_sc_hd__xor2_1 _0944_ (.A(_0339_),
    .B(_0386_),
    .X(_0468_));
 sky130_fd_sc_hd__o2111a_1 _0945_ (.A1(_0466_),
    .A2(_0467_),
    .B1(\dither.d_n_input[3] ),
    .C1(\dither.d_n_input[5] ),
    .D1(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_2 _0946_ (.A0(_0465_),
    .A1(_0463_),
    .S(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__o21a_1 _0947_ (.A1(_0363_),
    .A2(_0435_),
    .B1(_0444_),
    .X(\dither.d_n_input[7] ));
 sky130_fd_sc_hd__and3_1 _0948_ (.A(\dither.d_n_input[7] ),
    .B(_0469_),
    .C(_0463_),
    .X(_0471_));
 sky130_fd_sc_hd__a21oi_2 _0949_ (.A1(_0469_),
    .A2(_0463_),
    .B1(\dither.d_n_input[7] ),
    .Y(_0472_));
 sky130_fd_sc_hd__a211o_1 _0950_ (.A1(_0462_),
    .A2(_0470_),
    .B1(_0471_),
    .C1(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__o21a_1 _0951_ (.A1(_0385_),
    .A2(_0435_),
    .B1(_0444_),
    .X(\dither.d_n_input[8] ));
 sky130_fd_sc_hd__nor2_1 _0952_ (.A(_0471_),
    .B(\dither.d_n_input[8] ),
    .Y(_0474_));
 sky130_fd_sc_hd__or2_1 _0953_ (.A(_0473_),
    .B(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__inv_2 _0954_ (.A(\clkdivider.count[4] ),
    .Y(_0476_));
 sky130_fd_sc_hd__o211ai_2 _0955_ (.A1(_0471_),
    .A2(_0472_),
    .B1(_0462_),
    .C1(_0470_),
    .Y(_0477_));
 sky130_fd_sc_hd__and3_1 _0956_ (.A(_0476_),
    .B(_0473_),
    .C(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__inv_2 _0957_ (.A(\clkdivider.count[2] ),
    .Y(_0479_));
 sky130_fd_sc_hd__o21a_1 _0958_ (.A1(_0460_),
    .A2(\dither.d_n_input[4] ),
    .B1(_0461_),
    .X(_0480_));
 sky130_fd_sc_hd__xnor2_2 _0959_ (.A(_0461_),
    .B(\dither.d_n_input[5] ),
    .Y(_0481_));
 sky130_fd_sc_hd__o21a_1 _0960_ (.A1(_0480_),
    .A2(_0481_),
    .B1(_0462_),
    .X(_0482_));
 sky130_fd_sc_hd__a21o_1 _0961_ (.A1(_0451_),
    .A2(_0458_),
    .B1(_0459_),
    .X(_0483_));
 sky130_fd_sc_hd__inv_2 _0962_ (.A(net21),
    .Y(_0011_));
 sky130_fd_sc_hd__o31a_1 _0963_ (.A1(_0466_),
    .A2(_0467_),
    .A3(\dither.d_n_input[3] ),
    .B1(_0011_),
    .X(_0484_));
 sky130_fd_sc_hd__and3b_1 _0964_ (.A_N(\clkdivider.count[1] ),
    .B(_0483_),
    .C(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__or2b_1 _0965_ (.A(_0485_),
    .B_N(_0480_),
    .X(_0486_));
 sky130_fd_sc_hd__a21bo_1 _0966_ (.A1(_0483_),
    .A2(_0484_),
    .B1_N(\clkdivider.count[1] ),
    .X(_0487_));
 sky130_fd_sc_hd__o211a_1 _0967_ (.A1(_0479_),
    .A2(_0482_),
    .B1(_0486_),
    .C1(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__and2_1 _0968_ (.A(_0462_),
    .B(_0470_),
    .X(_0489_));
 sky130_fd_sc_hd__nor2_1 _0969_ (.A(_0462_),
    .B(_0470_),
    .Y(_0490_));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(\clkdivider.count[3] ),
    .Y(_0491_));
 sky130_fd_sc_hd__o21a_1 _0971_ (.A1(_0489_),
    .A2(_0490_),
    .B1(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__and2_1 _0972_ (.A(_0479_),
    .B(_0482_),
    .X(_0493_));
 sky130_fd_sc_hd__or3_1 _0973_ (.A(_0491_),
    .B(_0489_),
    .C(_0490_),
    .X(_0494_));
 sky130_fd_sc_hd__a21o_1 _0974_ (.A1(_0473_),
    .A2(_0477_),
    .B1(_0476_),
    .X(_0495_));
 sky130_fd_sc_hd__o311a_1 _0975_ (.A1(_0488_),
    .A2(_0492_),
    .A3(_0493_),
    .B1(_0494_),
    .C1(_0495_),
    .X(_0496_));
 sky130_fd_sc_hd__xnor2_1 _0976_ (.A(_0473_),
    .B(_0474_),
    .Y(_0497_));
 sky130_fd_sc_hd__a2bb2o_1 _0977_ (.A1_N(_0478_),
    .A2_N(_0496_),
    .B1(\clkdivider.count[5] ),
    .B2(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__o22a_1 _0978_ (.A1(\clkdivider.count[6] ),
    .A2(_0475_),
    .B1(_0497_),
    .B2(\clkdivider.count[5] ),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_1 _0979_ (.A(\clkdivider.count[5] ),
    .B(\clkdivider.count[6] ),
    .Y(_0500_));
 sky130_fd_sc_hd__or4_1 _0980_ (.A(\clkdivider.count[4] ),
    .B(\clkdivider.count[0] ),
    .C(\clkdivider.count[1] ),
    .D(\clkdivider.count[6] ),
    .X(_0501_));
 sky130_fd_sc_hd__or4_1 _0981_ (.A(\clkdivider.count[3] ),
    .B(\clkdivider.count[2] ),
    .C(\clkdivider.count[5] ),
    .D(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__o211a_1 _0982_ (.A1(_0476_),
    .A2(_0500_),
    .B1(_0502_),
    .C1(net34),
    .X(_0503_));
 sky130_fd_sc_hd__a221o_1 _0983_ (.A1(net26),
    .A2(_0475_),
    .B1(_0498_),
    .B2(_0499_),
    .C1(_0503_),
    .X(_0080_));
 sky130_fd_sc_hd__inv_2 _0984_ (.A(net11),
    .Y(_0504_));
 sky130_fd_sc_hd__nand2_1 _0985_ (.A(_0469_),
    .B(_0463_),
    .Y(_0505_));
 sky130_fd_sc_hd__o21a_1 _0986_ (.A1(_0469_),
    .A2(\dither.d_n_input[6] ),
    .B1(_0505_),
    .X(_0506_));
 sky130_fd_sc_hd__a221o_1 _0987_ (.A1(_0479_),
    .A2(_0481_),
    .B1(_0487_),
    .B2(_0480_),
    .C1(_0485_),
    .X(_0507_));
 sky130_fd_sc_hd__o221ai_2 _0988_ (.A1(_0491_),
    .A2(_0506_),
    .B1(_0481_),
    .B2(_0479_),
    .C1(_0507_),
    .Y(_0508_));
 sky130_fd_sc_hd__or2_1 _0989_ (.A(_0471_),
    .B(_0472_),
    .X(_0509_));
 sky130_fd_sc_hd__o22a_1 _0990_ (.A1(\clkdivider.count[4] ),
    .A2(_0509_),
    .B1(_0470_),
    .B2(\clkdivider.count[3] ),
    .X(_0510_));
 sky130_fd_sc_hd__a22o_1 _0991_ (.A1(\clkdivider.count[4] ),
    .A2(_0509_),
    .B1(_0474_),
    .B2(\clkdivider.count[5] ),
    .X(_0511_));
 sky130_fd_sc_hd__a21o_1 _0992_ (.A1(_0508_),
    .A2(_0510_),
    .B1(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__or2_1 _0993_ (.A(\clkdivider.count[5] ),
    .B(_0474_),
    .X(_0513_));
 sky130_fd_sc_hd__a221oi_1 _0994_ (.A1(_0504_),
    .A2(_0502_),
    .B1(_0512_),
    .B2(_0513_),
    .C1(net26),
    .Y(_0079_));
 sky130_fd_sc_hd__or4_1 _0995_ (.A(\clkdivider.count[3] ),
    .B(\clkdivider.count[2] ),
    .C(_0476_),
    .D(\clkdivider.count[5] ),
    .X(_0514_));
 sky130_fd_sc_hd__buf_1 _0996_ (.A(_0514_),
    .X(_0000_));
 sky130_fd_sc_hd__inv_2 _0997_ (.A(_0455_),
    .Y(\dither.d_n_input[2] ));
 sky130_fd_sc_hd__and4_1 _0998_ (.A(\clkdivider.count[3] ),
    .B(\clkdivider.count[2] ),
    .C(\clkdivider.count[4] ),
    .D(\clkdivider.count[5] ),
    .X(_0515_));
 sky130_fd_sc_hd__clkbuf_1 _0999_ (.A(_0515_),
    .X(_0007_));
 sky130_fd_sc_hd__nand2_1 _1000_ (.A(\dither.count[1] ),
    .B(\dither.count[0] ),
    .Y(_0516_));
 sky130_fd_sc_hd__or2_1 _1001_ (.A(\dither.count[1] ),
    .B(\dither.count[0] ),
    .X(_0517_));
 sky130_fd_sc_hd__and2_1 _1002_ (.A(_0516_),
    .B(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_1 _1003_ (.A(_0518_),
    .X(_0009_));
 sky130_fd_sc_hd__xnor2_1 _1004_ (.A(\dither.count[2] ),
    .B(_0516_),
    .Y(_0010_));
 sky130_fd_sc_hd__xor2_1 _1005_ (.A(net21),
    .B(net28),
    .X(_0012_));
 sky130_fd_sc_hd__and3_1 _1006_ (.A(\clkdivider.count[2] ),
    .B(\clkdivider.count[0] ),
    .C(\clkdivider.count[1] ),
    .X(_0519_));
 sky130_fd_sc_hd__a21oi_1 _1007_ (.A1(net21),
    .A2(net28),
    .B1(net32),
    .Y(_0520_));
 sky130_fd_sc_hd__nor2_1 _1008_ (.A(_0519_),
    .B(_0520_),
    .Y(_0013_));
 sky130_fd_sc_hd__nand2_1 _1009_ (.A(\clkdivider.count[3] ),
    .B(_0519_),
    .Y(_0521_));
 sky130_fd_sc_hd__or2_1 _1010_ (.A(\clkdivider.count[3] ),
    .B(_0519_),
    .X(_0522_));
 sky130_fd_sc_hd__and2_1 _1011_ (.A(_0521_),
    .B(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_1 _1012_ (.A(_0523_),
    .X(_0014_));
 sky130_fd_sc_hd__xnor2_1 _1013_ (.A(net33),
    .B(_0521_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand4_1 _1014_ (.A(\clkdivider.count[3] ),
    .B(\clkdivider.count[4] ),
    .C(\clkdivider.count[5] ),
    .D(_0519_),
    .Y(_0524_));
 sky130_fd_sc_hd__a31o_1 _1015_ (.A1(\clkdivider.count[3] ),
    .A2(\clkdivider.count[4] ),
    .A3(_0519_),
    .B1(\clkdivider.count[5] ),
    .X(_0525_));
 sky130_fd_sc_hd__and2_1 _1016_ (.A(_0524_),
    .B(_0525_),
    .X(_0526_));
 sky130_fd_sc_hd__clkbuf_1 _1017_ (.A(_0526_),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _1018_ (.A(\clkdivider.count[6] ),
    .B(_0524_),
    .X(_0527_));
 sky130_fd_sc_hd__clkbuf_1 _1019_ (.A(_0527_),
    .X(_0017_));
 sky130_fd_sc_hd__and2b_1 _1020_ (.A_N(_0173_),
    .B(_0172_),
    .X(_0528_));
 sky130_fd_sc_hd__xnor2_1 _1021_ (.A(_0170_),
    .B(_0528_),
    .Y(_0529_));
 sky130_fd_sc_hd__a21oi_1 _1022_ (.A1(_0450_),
    .A2(_0529_),
    .B1(_0445_),
    .Y(\stanley.d_n_reg[0] ));
 sky130_fd_sc_hd__nor2_1 _1023_ (.A(_0394_),
    .B(_0453_),
    .Y(\stanley.d_n_reg[1] ));
 sky130_fd_sc_hd__a21oi_1 _1024_ (.A1(_0393_),
    .A2(_0450_),
    .B1(_0445_),
    .Y(\stanley.d_n_reg[2] ));
 sky130_fd_sc_hd__nor2_1 _1025_ (.A(_0391_),
    .B(_0392_),
    .Y(_0530_));
 sky130_fd_sc_hd__o21a_1 _1026_ (.A1(_0530_),
    .A2(_0453_),
    .B1(_0444_),
    .X(\stanley.d_n_reg[3] ));
 sky130_fd_sc_hd__nor2_1 _1027_ (.A(_0397_),
    .B(_0453_),
    .Y(\stanley.d_n_reg[4] ));
 sky130_fd_sc_hd__nor2_1 _1028_ (.A(_0396_),
    .B(_0453_),
    .Y(\stanley.d_n_reg[5] ));
 sky130_fd_sc_hd__o21ai_1 _1029_ (.A1(net6),
    .A2(net5),
    .B1(net7),
    .Y(_0531_));
 sky130_fd_sc_hd__a21o_1 _1030_ (.A1(net6),
    .A2(net5),
    .B1(net7),
    .X(_0532_));
 sky130_fd_sc_hd__and3_1 _1031_ (.A(net8),
    .B(_0531_),
    .C(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__or3_1 _1032_ (.A(net2),
    .B(net1),
    .C(net3),
    .X(_0534_));
 sky130_fd_sc_hd__o21ai_1 _1033_ (.A1(net2),
    .A2(net1),
    .B1(net3),
    .Y(_0535_));
 sky130_fd_sc_hd__and3_1 _1034_ (.A(_0533_),
    .B(_0534_),
    .C(_0535_),
    .X(_0536_));
 sky130_fd_sc_hd__clkbuf_1 _1035_ (.A(_0536_),
    .X(_0018_));
 sky130_fd_sc_hd__or2_1 _1036_ (.A(net4),
    .B(_0534_),
    .X(_0537_));
 sky130_fd_sc_hd__nand2_1 _1037_ (.A(net4),
    .B(_0534_),
    .Y(_0538_));
 sky130_fd_sc_hd__and3_1 _1038_ (.A(_0533_),
    .B(_0537_),
    .C(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_1 _1039_ (.A(_0539_),
    .X(_0019_));
 sky130_fd_sc_hd__o311a_1 _1040_ (.A1(net6),
    .A2(net5),
    .A3(_0537_),
    .B1(net7),
    .C1(net8),
    .X(_0021_));
 sky130_fd_sc_hd__a31o_1 _1041_ (.A1(net6),
    .A2(net5),
    .A3(_0537_),
    .B1(net7),
    .X(_0540_));
 sky130_fd_sc_hd__nand3b_1 _1042_ (.A_N(_0021_),
    .B(net8),
    .C(_0540_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _1043_ (.A(net20),
    .Y(_0001_));
 sky130_fd_sc_hd__xor2_1 _1044_ (.A(net24),
    .B(net20),
    .X(_0002_));
 sky130_fd_sc_hd__a21oi_1 _1045_ (.A1(\clkdivider.clk2[1] ),
    .A2(\clkdivider.clk2[0] ),
    .B1(net22),
    .Y(_0541_));
 sky130_fd_sc_hd__nor2_1 _1046_ (.A(_0082_),
    .B(net23),
    .Y(_0003_));
 sky130_fd_sc_hd__nor2_1 _1047_ (.A(net25),
    .B(_0082_),
    .Y(_0542_));
 sky130_fd_sc_hd__nor2_1 _1048_ (.A(_0083_),
    .B(_0542_),
    .Y(_0004_));
 sky130_fd_sc_hd__xor2_1 _1049_ (.A(net19),
    .B(_0083_),
    .X(_0005_));
 sky130_fd_sc_hd__and2_1 _1050_ (.A(net31),
    .B(_0084_),
    .X(_0543_));
 sky130_fd_sc_hd__clkbuf_1 _1051_ (.A(_0543_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_4 _1052_ (.A(net9),
    .X(_0544_));
 sky130_fd_sc_hd__buf_4 _1053_ (.A(_0544_),
    .X(_0545_));
 sky130_fd_sc_hd__inv_2 _1054_ (.A(_0545_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1055_ (.A(_0545_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1056_ (.A(_0545_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1057_ (.A(_0545_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1058_ (.A(_0545_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1059_ (.A(_0545_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1060_ (.A(_0545_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1061_ (.A(_0545_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1062_ (.A(_0545_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _1063_ (.A(_0545_),
    .Y(_0031_));
 sky130_fd_sc_hd__clkbuf_8 _1064_ (.A(_0544_),
    .X(_0546_));
 sky130_fd_sc_hd__inv_2 _1065_ (.A(_0546_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1066_ (.A(_0546_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1067_ (.A(_0546_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(_0546_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(_0546_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1070_ (.A(_0546_),
    .Y(_0037_));
 sky130_fd_sc_hd__inv_2 _1071_ (.A(_0546_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1072_ (.A(_0546_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(_0546_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1074_ (.A(_0546_),
    .Y(_0041_));
 sky130_fd_sc_hd__clkbuf_8 _1075_ (.A(_0544_),
    .X(_0547_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(_0547_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(_0547_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1078_ (.A(_0547_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1079_ (.A(_0547_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1080_ (.A(_0547_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1081_ (.A(_0547_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1082_ (.A(_0547_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1083_ (.A(_0547_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _1084_ (.A(_0547_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _1085_ (.A(_0547_),
    .Y(_0051_));
 sky130_fd_sc_hd__buf_4 _1086_ (.A(net9),
    .X(_0548_));
 sky130_fd_sc_hd__inv_2 _1087_ (.A(_0548_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _1088_ (.A(_0548_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _1089_ (.A(_0548_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _1090_ (.A(_0548_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _1091_ (.A(_0548_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _1092_ (.A(_0548_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _1093_ (.A(_0548_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _1094_ (.A(_0548_),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _1095_ (.A(_0548_),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _1096_ (.A(_0548_),
    .Y(_0061_));
 sky130_fd_sc_hd__buf_4 _1097_ (.A(net9),
    .X(_0549_));
 sky130_fd_sc_hd__inv_2 _1098_ (.A(_0549_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _1099_ (.A(_0549_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _1100_ (.A(_0549_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _1101_ (.A(_0549_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _1102_ (.A(_0549_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _1103_ (.A(_0549_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _1104_ (.A(_0549_),
    .Y(_0068_));
 sky130_fd_sc_hd__inv_2 _1105_ (.A(_0549_),
    .Y(_0069_));
 sky130_fd_sc_hd__inv_2 _1106_ (.A(_0549_),
    .Y(_0070_));
 sky130_fd_sc_hd__inv_2 _1107_ (.A(_0549_),
    .Y(_0071_));
 sky130_fd_sc_hd__inv_2 _1108_ (.A(_0544_),
    .Y(_0072_));
 sky130_fd_sc_hd__inv_2 _1109_ (.A(_0544_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _1110_ (.A(_0544_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1111_ (.A(_0544_),
    .Y(_0075_));
 sky130_fd_sc_hd__inv_2 _1112_ (.A(_0544_),
    .Y(_0076_));
 sky130_fd_sc_hd__inv_2 _1113_ (.A(_0544_),
    .Y(_0077_));
 sky130_fd_sc_hd__inv_2 _1114_ (.A(_0544_),
    .Y(_0078_));
 sky130_fd_sc_hd__dfrtp_1 _1115_ (.CLK(clknet_1_1__leaf_clk),
    .D(net27),
    .RESET_B(_0022_),
    .Q(net11));
 sky130_fd_sc_hd__dfrtp_4 _1116_ (.CLK(\clkdivider.clk_dpwm ),
    .D(_0008_),
    .RESET_B(_0023_),
    .Q(\dither.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1117_ (.CLK(\clkdivider.clk_dpwm ),
    .D(_0009_),
    .RESET_B(_0024_),
    .Q(\dither.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1118_ (.CLK(\clkdivider.clk_dpwm ),
    .D(_0010_),
    .RESET_B(_0025_),
    .Q(\dither.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1119_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0011_),
    .RESET_B(_0026_),
    .Q(\clkdivider.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1120_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0012_),
    .RESET_B(_0027_),
    .Q(\clkdivider.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _1121_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0013_),
    .RESET_B(_0028_),
    .Q(\clkdivider.count[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1122_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0014_),
    .RESET_B(_0029_),
    .Q(\clkdivider.count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1123_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0015_),
    .RESET_B(_0030_),
    .Q(\clkdivider.count[4] ));
 sky130_fd_sc_hd__dfrtp_4 _1124_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0016_),
    .RESET_B(_0031_),
    .Q(\clkdivider.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1125_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0017_),
    .RESET_B(_0032_),
    .Q(\clkdivider.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1126_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0080_),
    .RESET_B(_0033_),
    .Q(net12));
 sky130_fd_sc_hd__dfrtp_1 _1127_ (.CLK(clknet_1_1__leaf_clk),
    .D(net30),
    .RESET_B(_0034_),
    .Q(\clkdivider.clk_dpwm ));
 sky130_fd_sc_hd__dfrtp_1 _1128_ (.CLK(net17),
    .D(\stanley.d_n_reg[0] ),
    .RESET_B(_0035_),
    .Q(\stanley.d_n_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1129_ (.CLK(net17),
    .D(\stanley.d_n_reg[1] ),
    .RESET_B(_0036_),
    .Q(\stanley.d_n_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1130_ (.CLK(net17),
    .D(\stanley.d_n_reg[2] ),
    .RESET_B(_0037_),
    .Q(\stanley.d_n_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1131_ (.CLK(net17),
    .D(\stanley.d_n_reg[3] ),
    .RESET_B(_0038_),
    .Q(\stanley.d_n_1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1132_ (.CLK(net17),
    .D(\stanley.d_n_reg[4] ),
    .RESET_B(_0039_),
    .Q(\stanley.d_n_1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1133_ (.CLK(net17),
    .D(\stanley.d_n_reg[5] ),
    .RESET_B(_0040_),
    .Q(\stanley.d_n_1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1134_ (.CLK(net16),
    .D(\dither.d_n_input[0] ),
    .RESET_B(_0041_),
    .Q(\stanley.d_n_1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1135_ (.CLK(net16),
    .D(\dither.d_n_input[1] ),
    .RESET_B(_0042_),
    .Q(\stanley.d_n_1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1136_ (.CLK(net16),
    .D(\dither.d_n_input[2] ),
    .RESET_B(_0043_),
    .Q(\stanley.d_n_1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _1137_ (.CLK(net16),
    .D(\dither.d_n_input[3] ),
    .RESET_B(_0044_),
    .Q(\stanley.d_n_1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _1138_ (.CLK(net16),
    .D(\dither.d_n_input[4] ),
    .RESET_B(_0045_),
    .Q(\stanley.d_n_1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _1139_ (.CLK(net16),
    .D(\dither.d_n_input[5] ),
    .RESET_B(_0046_),
    .Q(\stanley.d_n_1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _1140_ (.CLK(net16),
    .D(\dither.d_n_input[6] ),
    .RESET_B(_0047_),
    .Q(\stanley.d_n_1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1141_ (.CLK(net16),
    .D(\dither.d_n_input[7] ),
    .RESET_B(_0048_),
    .Q(\stanley.d_n_1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1142_ (.CLK(net16),
    .D(\dither.d_n_input[8] ),
    .RESET_B(_0049_),
    .Q(\stanley.d_n_1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1143_ (.CLK(net16),
    .D(net18),
    .RESET_B(_0050_),
    .Q(\stanley.d_n_1[15] ));
 sky130_fd_sc_hd__conb_1 _1143__18 (.LO(net18));
 sky130_fd_sc_hd__dfrtp_4 _1144_ (.CLK(net17),
    .D(\stanley.en2[0] ),
    .RESET_B(_0051_),
    .Q(\stanley.en3[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1145_ (.CLK(net14),
    .D(\stanley.en2[1] ),
    .RESET_B(_0052_),
    .Q(\stanley.en3[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1146_ (.CLK(net14),
    .D(\stanley.en2[2] ),
    .RESET_B(_0053_),
    .Q(\stanley.en3[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1147_ (.CLK(net15),
    .D(\stanley.en2[3] ),
    .RESET_B(_0054_),
    .Q(\stanley.en3[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1148_ (.CLK(net14),
    .D(\stanley.en1[0] ),
    .RESET_B(_0055_),
    .Q(\stanley.en2[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1149_ (.CLK(net14),
    .D(\stanley.en1[1] ),
    .RESET_B(_0056_),
    .Q(\stanley.en2[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1150_ (.CLK(net14),
    .D(\stanley.en1[2] ),
    .RESET_B(_0057_),
    .Q(\stanley.en2[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1151_ (.CLK(net14),
    .D(net13),
    .RESET_B(_0058_),
    .Q(\stanley.en2[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1152_ (.CLK(net14),
    .D(\stanley.en[0] ),
    .RESET_B(_0059_),
    .Q(\stanley.en1[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1153_ (.CLK(net14),
    .D(\stanley.en[1] ),
    .RESET_B(_0060_),
    .Q(\stanley.en1[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1154_ (.CLK(net14),
    .D(\stanley.en[2] ),
    .RESET_B(_0061_),
    .Q(\stanley.en1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1155_ (.CLK(net14),
    .D(\stanley.en[3] ),
    .RESET_B(_0062_),
    .Q(\stanley.en1[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1156_ (.CLK(net15),
    .D(\encoder.en[0] ),
    .RESET_B(_0063_),
    .Q(\stanley.en[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1157_ (.CLK(net15),
    .D(\encoder.en[1] ),
    .RESET_B(_0064_),
    .Q(\stanley.en[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1158_ (.CLK(net15),
    .D(\encoder.en[2] ),
    .RESET_B(_0065_),
    .Q(\stanley.en[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1159_ (.CLK(net15),
    .D(\encoder.en[3] ),
    .RESET_B(_0066_),
    .Q(\stanley.en[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1160_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0018_),
    .RESET_B(_0067_),
    .Q(\encoder.en[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1161_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0019_),
    .RESET_B(_0068_),
    .Q(\encoder.en[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1162_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0020_),
    .RESET_B(_0069_),
    .Q(\encoder.en[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1163_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0021_),
    .RESET_B(_0070_),
    .Q(\encoder.en[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1164_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0000_),
    .RESET_B(_0071_),
    .Q(net10));
 sky130_fd_sc_hd__dfrtp_4 _1165_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0007_),
    .RESET_B(_0072_),
    .Q(\clkdivider.clk_comp ));
 sky130_fd_sc_hd__dfrtp_1 _1166_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0001_),
    .RESET_B(_0073_),
    .Q(\clkdivider.clk2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1167_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0002_),
    .RESET_B(_0074_),
    .Q(\clkdivider.clk2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1168_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0003_),
    .RESET_B(_0075_),
    .Q(\clkdivider.clk2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1169_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0004_),
    .RESET_B(_0076_),
    .Q(\clkdivider.clk2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1170_ (.CLK(clknet_1_1__leaf_clk),
    .D(_0005_),
    .RESET_B(_0077_),
    .Q(\clkdivider.clk2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1171_ (.CLK(clknet_1_0__leaf_clk),
    .D(_0006_),
    .RESET_B(_0078_),
    .Q(\clkdivider.clk2[5] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_clk (.A(clknet_0_clk),
    .X(clknet_1_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_clk (.A(clknet_0_clk),
    .X(clknet_1_1__leaf_clk));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(\stanley.en1[3] ),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(net15),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(\clkdivider.clk_comp ),
    .X(net15));
 sky130_fd_sc_hd__buf_2 fanout16 (.A(\clkdivider.clk_comp ),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 fanout17 (.A(\clkdivider.clk_comp ),
    .X(net17));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\clkdivider.clk2[4] ),
    .X(net19));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\clkdivider.count[1] ),
    .X(net28));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\clkdivider.clk_dpwm ),
    .X(net29));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0081_),
    .X(net30));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\clkdivider.clk2[5] ),
    .X(net31));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\clkdivider.count[2] ),
    .X(net32));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\clkdivider.count[4] ),
    .X(net33));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net12),
    .X(net34));
 sky130_fd_sc_hd__buf_1 hold2 (.A(\clkdivider.clk2[0] ),
    .X(net20));
 sky130_fd_sc_hd__buf_1 hold3 (.A(\clkdivider.count[0] ),
    .X(net21));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\clkdivider.clk2[2] ),
    .X(net22));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0541_),
    .X(net23));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\clkdivider.clk2[1] ),
    .X(net24));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\clkdivider.clk2[3] ),
    .X(net25));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\clkdivider.count[6] ),
    .X(net26));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0079_),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(data_in[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(data_in[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(data_in[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(data_in[3]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(data_in[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(data_in[5]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(data_in[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(data_in[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(rst),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 output10 (.A(net10),
    .X(convst_bar));
 sky130_fd_sc_hd__clkbuf_4 output11 (.A(net11),
    .X(duty_high));
 sky130_fd_sc_hd__clkbuf_4 output12 (.A(net12),
    .X(duty_low));
endmodule

