library verilog;
use verilog.vl_types.all;
entity dither is
    port(
        clk_in          : in     vl_logic;
        rst             : in     vl_logic;
        d_n_input       : in     vl_logic_vector(8 downto 0);
        d_dith          : out    vl_logic_vector(5 downto 0)
    );
end dither;
